`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
module Fulladder1bit(
    input A, B, Cin,
    output Z, Cout
    );

assign Z= A^B^Cin;
assign Cout = A&B | B&Cin | Cin&A;


endmodule
